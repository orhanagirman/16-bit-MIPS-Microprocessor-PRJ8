----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:42:57 08/28/2020 
-- Design Name: 
-- Module Name:    pc - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity data_memory is
    Port ( clk : in  STD_LOGIC;
	        rst : in  STD_LOGIC;
			  dd : in  STD_LOGIC_VECTOR (15 downto 0);
			  mWrite : in STD_LOGIC;
           read_data : out  STD_LOGIC_VECTOR (15 downto 0));
end data_memory;

architecture Behavioral of data_memory is

begin
     process(clk,rst)
	  begin
	       if (rst = '1') then 
			     read_data <= "0000000000000000";
			 else
			     if (mWrite = '1') then
                  if rising_edge(clk) then
					      read_data <= dd;
				      end if;
              end if;						
          end if;
    end process;
end Behavioral;
